/*
 * DE0Nano_Button.v
 *
 *  ___       _         _   _       _ ___ _ _ ___
 *	| __._ _ _| |_ ___ _| |_| |___ _| | . | \ |_ _|
 *	| _>| ' ' | . / ._/ . / . / ._/ . |   |   || |
 *	|___|_|_|_|___\___\___\___\___\___|_|_|_\_||_|
 *
 *
 *  Created on	: 20/06/2015
 *      Author	: Ernesto Andres Rincon Cruz
 *      Web		: www.embeddedant.org
 *		  Device : EP4CE22F17C6N
 *		  Board  : DEO-NANO
 *
 *      Revision History:
 *			Rev 1.0.0 - (ErnestoARC) First release 20/06/2015.
 */ 
//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE0Nano_Button(
	//////////// CLOCK //////////
	CLOCK_50,
	//////////// LED //////////
	LED,
	//////////// KEY //////////
	KEY 
);

//=======================================================
//  PARAMETER declarations
//=======================================================
parameter LED_SEQUENCE_0		=8'b10000000;	
parameter LED_SEQUENCE_1		=8'b01000000;	
parameter LED_SEQUENCE_2		=8'b00100000;	
parameter LED_SEQUENCE_3		=8'b00010000;	
parameter LED_SEQUENCE_4		=8'b00001000;	
parameter LED_SEQUENCE_5		=8'b00000100;	
parameter LED_SEQUENCE_6		=8'b00000010;	
parameter LED_SEQUENCE_7		=8'b00000001;	

//=======================================================
//  PORT declarations
//=======================================================
//////////// CLOCK //////////
input 		          		CLOCK_50;
//////////// LED //////////
output		     [7:0]		LED;
//////////// KEY //////////
input 		     [1:0]		KEY;

//=======================================================
//  REG/WIRE declarations
//=======================================================
reg	[7:0]LedsState=LED_SEQUENCE_0;
reg	[7:0]LedsNextState;
wire 	Clock_Sequence;

reg	SequenceControl=0;
wire  Btn1_Signal;
wire  Btn2_Signal;


//Frequency Divider Module
ClockDivider #(.Bits_counter (28)) DIVIDER_A
	 (	.P_CLOCK(CLOCK_50),
		.P_TIMER_OUT(Clock_Sequence),
		.P_COMPARATOR(28'd16000000));
		
// Debounce circuir for Button1		
 DeBounce DebBtn1 (
        .clk(CLOCK_50), 
        .n_reset(1'b1), 
        .button_in(KEY[0]), 
        .DB_out(Btn1_Signal)
        );
		  
// Debounce circuir for Button2	  
 DeBounce DebBtn2 (
        .clk(CLOCK_50), 
        .n_reset(1'b1), 
        .button_in(KEY[1]), 
        .DB_out(Btn2_Signal)
        );  
//=======================================================
//  Structural coding
//=======================================================

	// Leds Sequence control 
	always @(*)
	begin
		case (LedsState)	
			LED_SEQUENCE_0:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_1;
					else	
						LedsNextState=LED_SEQUENCE_7;
				end
					
			LED_SEQUENCE_1:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_2;
					else	
						LedsNextState=LED_SEQUENCE_0;
				end

			LED_SEQUENCE_2:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_3;
					else	
						LedsNextState=LED_SEQUENCE_1;
				end
				
			LED_SEQUENCE_3:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_4;
					else	
						LedsNextState=LED_SEQUENCE_2;
				end
				
			LED_SEQUENCE_4:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_5;
					else	
						LedsNextState=LED_SEQUENCE_3;
				end
				
			LED_SEQUENCE_5:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_6;
					else	
						LedsNextState=LED_SEQUENCE_4;
				end
				
			LED_SEQUENCE_6:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_7;
					else	
						LedsNextState=LED_SEQUENCE_5;
				end
				
			LED_SEQUENCE_7:
				begin
					if (SequenceControl==0)
						LedsNextState=LED_SEQUENCE_0;
					else	
						LedsNextState=LED_SEQUENCE_6;
				end
				
			default:
						LedsNextState=LED_SEQUENCE_0;
		endcase
	end
	
	
	// Led direction control
	always @ (posedge CLOCK_50)
	begin
		if (Btn1_Signal==0)
			SequenceControl<=0;
		else if 	(Btn2_Signal==0)
			SequenceControl<=1;
		else 	
			SequenceControl<=SequenceControl;
	end
	
	
	// Leds sequence registers
	always @ (posedge Clock_Sequence)
	begin
		LedsState<=LedsNextState;
	end
//=======================================================
// 			Connections & assigns
//=======================================================
assign	LED 	= LedsState;

endmodule
