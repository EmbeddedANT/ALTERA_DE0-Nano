/*
 * DE0-Nano_Leds.v
 *
 *  ___       _         _   _       _ ___ _ _ ___
 *	| __._ _ _| |_ ___ _| |_| |___ _| | . | \ |_ _|
 *	| _>| ' ' | . / ._/ . / . / ._/ . |   |   || |
 *	|___|_|_|_|___\___\___\___\___\___|_|_|_\_||_|
 *
 *
 *  Created on	: 19/06/2015
 *      Author	: Ernesto Andres Rincon Cruz
 *      Web		: www.embeddedant.org
 *		  Device : EP4CE22F17C6N
 *		  Board  : DEO-NANO
 *
 *      Revision History:
 *			Rev 1.0.0 - (ErnestoARC) First created 19/06/2015.
 */    
//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE0Nano_Leds(
	//////////// CLOCK //////////
	CLOCK_50,
	//////////// LED //////////
	LED 
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK //////////
input	CLOCK_50;

//////////// LED //////////
output	[7:0]LED;


//=======================================================
//  REG/WIRE declarations
//=======================================================
wire Clock_2Hz;
reg [7:0]Counter=8'h00;

//Frequency Divider 50MHz -> 1Hz
ClockDivider #(.Bits_counter (28)) unit8
	 (	.P_CLOCK(CLOCK_50),
		.P_TIMER_OUT(Clock_2Hz),
		.P_COMPARATOR(28'd25000000));
		
//=======================================================
//  Structural coding
//=======================================================

	/*Counter for Leds*/
	always @ (posedge Clock_2Hz) begin
		Counter<=Counter+1;
	end
	
//=======================================================
// 			Connections & assigns
//=======================================================
assign	LED 	= Counter;

endmodule
