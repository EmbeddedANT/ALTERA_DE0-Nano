/*
 * ClockDivider.v
 *
 *  ___       _         _   _       _ ___ _ _ ___
 *	| __._ _ _| |_ ___ _| |_| |___ _| | . | \ |_ _|
 *	| _>| ' ' | . / ._/ . / . / ._/ . |   |   || |
 *	|___|_|_|_|___\___\___\___\___\___|_|_|_\_||_|
 *
 *
 *  Created on	: 20/06/2015
 *      Author	: Ernesto Andres Rincon Cruz
 *      Web		: www.embeddedant.org
 *		  Device : EP4CE22F17C6N
 *		  Board  : DEO-NANO
 *
 *      Revision History:
 *			Rev 1.0.0 - (ErnestoARC) First release 20/06/2015.
 */    
//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE0Nano_Switch(
	//////////// CLOCK //////////
	CLOCK_50,
	//////////// LED //////////
	LED,
	//////////// SW //////////
	SW 
);

//=======================================================
//  PARAMETER declarations
//=======================================================
parameter LED_SEQUENCE_0		=11'b10000001_000;	
parameter LED_SEQUENCE_1		=11'b01000010_001;	
parameter LED_SEQUENCE_2		=11'b00100100_010;	
parameter LED_SEQUENCE_3		=11'b00011000_011;	
parameter LED_SEQUENCE_4		=11'b00100100_100;	
parameter LED_SEQUENCE_5		=11'b01000010_101;	
//=======================================================
//  PORT declarations
//=======================================================
//////////// CLOCK //////////
input		CLOCK_50;
//////////// LED //////////
output	[7:0]LED;
//////////// SW //////////
input		[3:0]SW;
//=======================================================
//  REG/WIRE declarations
//=======================================================
wire 	Clock_Sequence;
reg	[10:0]LedsState;
reg	[10:0]LedsNextState;
reg 	[27:0]ClockSetup;

//Frequency Divider Module
ClockDivider #(.Bits_counter (28)) unit8
	 (	.P_CLOCK(CLOCK_50),
		.P_TIMER_OUT(Clock_Sequence),
		.P_COMPARATOR(ClockSetup));
//=======================================================
//  Structural coding
//=======================================================
	
	// Time Control with Switch
	always @(*)
	begin
		case (SW)
			4'h0: ClockSetup = 28'd1000000;	//50M/1M -> 	50.0Hz 
			4'h1: ClockSetup = 28'd2000000;	//50M/2M -> 	25.0Hz
			4'h2: ClockSetup = 28'd3000000;	//50M/3M -> 	16.66Hz
			4'h3: ClockSetup = 28'd4000000;	//50M/4M -> 	12.5Hz
			4'h4: ClockSetup = 28'd5000000;	//50M/5M -> 	10.0Hz
			4'h5: ClockSetup = 28'd6000000;	//50M/6M -> 	8.33Hz
			4'h6: ClockSetup = 28'd7000000;	//50M/7M -> 	7.14Hz
			4'h7: ClockSetup = 28'd8000000;	//50M/8M -> 	6.25Hz
			4'h8: ClockSetup = 28'd9000000;	//50M/9M -> 	5.55Hz
			4'h9: ClockSetup = 28'd10000000;	//50M/10M -> 	5.00Hz
			4'hA: ClockSetup = 28'd11000000;	//50M/11M -> 	4.54Hz
			4'hB: ClockSetup = 28'd12000000;	//50M/12M -> 	4.16Hz
			4'hC: ClockSetup = 28'd13000000;	//50M/13M -> 	3.84Hz
			4'hD: ClockSetup = 28'd14000000;	//50M/14M -> 	3.57Hz
			4'hE: ClockSetup = 28'd15000000;	//50M/15M -> 	3.33Hz
			4'hF: ClockSetup = 28'd16000000;	//50M/16M -> 	3.12Hz
		endcase	
	end

	// Leds Sequence control 
	always @(*)
	begin
		case (LedsState)	
			LED_SEQUENCE_0:  LedsNextState=LED_SEQUENCE_1;
			LED_SEQUENCE_1:  LedsNextState=LED_SEQUENCE_2;
			LED_SEQUENCE_2:  LedsNextState=LED_SEQUENCE_3;
			LED_SEQUENCE_3:  LedsNextState=LED_SEQUENCE_4;
			LED_SEQUENCE_4:  LedsNextState=LED_SEQUENCE_5;
			LED_SEQUENCE_5:  LedsNextState=LED_SEQUENCE_0;	
		endcase
	end
	
	// Leds sequence registers
	always @ (posedge Clock_Sequence)
	begin
		LedsState<=LedsNextState;
	end
	
	
	
//=======================================================
// 			Connections & assigns
//=======================================================
assign	LED 	= LedsState[10:3];

endmodule
