/*
 * ClockDivider.v
 *
 *  ___       _         _   _       _ ___ _ _ ___
 *	| __._ _ _| |_ ___ _| |_| |___ _| | . | \ |_ _|
 *	| _>| ' ' | . / ._/ . / . / ._/ . |   |   || |
 *	|___|_|_|_|___\___\___\___\___\___|_|_|_\_||_|
 *
 *
 *  Created on	: 19/06/2015
 *      Author	: Ernesto Andres Rincon Cruz
 *      Web		: www.embeddedant.org
 *		  Device : EP4CE22F17C6N
 *		  Board  : DEO-NANO
 *
 *      Revision History:
 *			Rev 1.0.0 - (ErnestoARC) First created 19/06/2015.
 */    
module ClockDivider
	#(parameter Bits_counter = 32)
	 (	input  P_CLOCK,
		output P_TIMER_OUT,
		input  [Bits_counter-1:0] P_COMPARATOR);
//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================


//=======================================================
//  REG/WIRE declarations
//=======================================================
   reg [Bits_counter-1:0] r_Timer;
   reg r_Result;
	
//=======================================================
//  Structural coding
//=======================================================
   always @(posedge P_CLOCK)
	begin
		if (r_Timer >= P_COMPARATOR)
			begin
			     r_Result <= !r_Result;
			     r_Timer <= 0;
			end		
		else
		   begin
			     r_Timer <= r_Timer+1; 
				  r_Result <= r_Result;
		   end
	end	
//=======================================================
// 			Connections & assigns
//=======================================================
assign P_TIMER_OUT = r_Result; 

endmodule
